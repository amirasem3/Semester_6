SHIFT4L_inst : SHIFT4L PORT MAP (
		result	 => result_sig
	);
