pushbyte_inst : pushbyte PORT MAP (
		result	 => result_sig
	);
