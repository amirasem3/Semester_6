IOR_inst : IOR PORT MAP (
		result	 => result_sig
	);
