WIDE_inst : WIDE PORT MAP (
		result	 => result_sig
	);
