ZERO19BIT_inst : ZERO19BIT PORT MAP (
		result	 => result_sig
	);
