B_inst : B PORT MAP (
		result	 => result_sig
	);
