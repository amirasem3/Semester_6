NOP_inst : NOP PORT MAP (
		result	 => result_sig
	);
