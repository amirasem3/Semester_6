GOTO_inst : GOTO PORT MAP (
		result	 => result_sig
	);
