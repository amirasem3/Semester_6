LDC_W_inst : LDC_W PORT MAP (
		result	 => result_sig
	);
