IF_ICM_inst : IF_ICM PORT MAP (
		result	 => result_sig
	);
