DUP_inst : DUP PORT MAP (
		result	 => result_sig
	);
