-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: mux3to8_32bit.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.1.1 Build 189 12/02/2015 SJ Lite Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux3to8_32bit IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END mux3to8_32bit;


ARCHITECTURE SYN OF mux3to8_32bit IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (7 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
	sub_wire8    <= data0x(31 DOWNTO 0);
	sub_wire7    <= data1x(31 DOWNTO 0);
	sub_wire6    <= data2x(31 DOWNTO 0);
	sub_wire5    <= data3x(31 DOWNTO 0);
	sub_wire4    <= data4x(31 DOWNTO 0);
	sub_wire3    <= data5x(31 DOWNTO 0);
	sub_wire2    <= data6x(31 DOWNTO 0);
	sub_wire0    <= data7x(31 DOWNTO 0);
	sub_wire1(7, 0)    <= sub_wire0(0);
	sub_wire1(7, 1)    <= sub_wire0(1);
	sub_wire1(7, 2)    <= sub_wire0(2);
	sub_wire1(7, 3)    <= sub_wire0(3);
	sub_wire1(7, 4)    <= sub_wire0(4);
	sub_wire1(7, 5)    <= sub_wire0(5);
	sub_wire1(7, 6)    <= sub_wire0(6);
	sub_wire1(7, 7)    <= sub_wire0(7);
	sub_wire1(7, 8)    <= sub_wire0(8);
	sub_wire1(7, 9)    <= sub_wire0(9);
	sub_wire1(7, 10)    <= sub_wire0(10);
	sub_wire1(7, 11)    <= sub_wire0(11);
	sub_wire1(7, 12)    <= sub_wire0(12);
	sub_wire1(7, 13)    <= sub_wire0(13);
	sub_wire1(7, 14)    <= sub_wire0(14);
	sub_wire1(7, 15)    <= sub_wire0(15);
	sub_wire1(7, 16)    <= sub_wire0(16);
	sub_wire1(7, 17)    <= sub_wire0(17);
	sub_wire1(7, 18)    <= sub_wire0(18);
	sub_wire1(7, 19)    <= sub_wire0(19);
	sub_wire1(7, 20)    <= sub_wire0(20);
	sub_wire1(7, 21)    <= sub_wire0(21);
	sub_wire1(7, 22)    <= sub_wire0(22);
	sub_wire1(7, 23)    <= sub_wire0(23);
	sub_wire1(7, 24)    <= sub_wire0(24);
	sub_wire1(7, 25)    <= sub_wire0(25);
	sub_wire1(7, 26)    <= sub_wire0(26);
	sub_wire1(7, 27)    <= sub_wire0(27);
	sub_wire1(7, 28)    <= sub_wire0(28);
	sub_wire1(7, 29)    <= sub_wire0(29);
	sub_wire1(7, 30)    <= sub_wire0(30);
	sub_wire1(7, 31)    <= sub_wire0(31);
	sub_wire1(6, 0)    <= sub_wire2(0);
	sub_wire1(6, 1)    <= sub_wire2(1);
	sub_wire1(6, 2)    <= sub_wire2(2);
	sub_wire1(6, 3)    <= sub_wire2(3);
	sub_wire1(6, 4)    <= sub_wire2(4);
	sub_wire1(6, 5)    <= sub_wire2(5);
	sub_wire1(6, 6)    <= sub_wire2(6);
	sub_wire1(6, 7)    <= sub_wire2(7);
	sub_wire1(6, 8)    <= sub_wire2(8);
	sub_wire1(6, 9)    <= sub_wire2(9);
	sub_wire1(6, 10)    <= sub_wire2(10);
	sub_wire1(6, 11)    <= sub_wire2(11);
	sub_wire1(6, 12)    <= sub_wire2(12);
	sub_wire1(6, 13)    <= sub_wire2(13);
	sub_wire1(6, 14)    <= sub_wire2(14);
	sub_wire1(6, 15)    <= sub_wire2(15);
	sub_wire1(6, 16)    <= sub_wire2(16);
	sub_wire1(6, 17)    <= sub_wire2(17);
	sub_wire1(6, 18)    <= sub_wire2(18);
	sub_wire1(6, 19)    <= sub_wire2(19);
	sub_wire1(6, 20)    <= sub_wire2(20);
	sub_wire1(6, 21)    <= sub_wire2(21);
	sub_wire1(6, 22)    <= sub_wire2(22);
	sub_wire1(6, 23)    <= sub_wire2(23);
	sub_wire1(6, 24)    <= sub_wire2(24);
	sub_wire1(6, 25)    <= sub_wire2(25);
	sub_wire1(6, 26)    <= sub_wire2(26);
	sub_wire1(6, 27)    <= sub_wire2(27);
	sub_wire1(6, 28)    <= sub_wire2(28);
	sub_wire1(6, 29)    <= sub_wire2(29);
	sub_wire1(6, 30)    <= sub_wire2(30);
	sub_wire1(6, 31)    <= sub_wire2(31);
	sub_wire1(5, 0)    <= sub_wire3(0);
	sub_wire1(5, 1)    <= sub_wire3(1);
	sub_wire1(5, 2)    <= sub_wire3(2);
	sub_wire1(5, 3)    <= sub_wire3(3);
	sub_wire1(5, 4)    <= sub_wire3(4);
	sub_wire1(5, 5)    <= sub_wire3(5);
	sub_wire1(5, 6)    <= sub_wire3(6);
	sub_wire1(5, 7)    <= sub_wire3(7);
	sub_wire1(5, 8)    <= sub_wire3(8);
	sub_wire1(5, 9)    <= sub_wire3(9);
	sub_wire1(5, 10)    <= sub_wire3(10);
	sub_wire1(5, 11)    <= sub_wire3(11);
	sub_wire1(5, 12)    <= sub_wire3(12);
	sub_wire1(5, 13)    <= sub_wire3(13);
	sub_wire1(5, 14)    <= sub_wire3(14);
	sub_wire1(5, 15)    <= sub_wire3(15);
	sub_wire1(5, 16)    <= sub_wire3(16);
	sub_wire1(5, 17)    <= sub_wire3(17);
	sub_wire1(5, 18)    <= sub_wire3(18);
	sub_wire1(5, 19)    <= sub_wire3(19);
	sub_wire1(5, 20)    <= sub_wire3(20);
	sub_wire1(5, 21)    <= sub_wire3(21);
	sub_wire1(5, 22)    <= sub_wire3(22);
	sub_wire1(5, 23)    <= sub_wire3(23);
	sub_wire1(5, 24)    <= sub_wire3(24);
	sub_wire1(5, 25)    <= sub_wire3(25);
	sub_wire1(5, 26)    <= sub_wire3(26);
	sub_wire1(5, 27)    <= sub_wire3(27);
	sub_wire1(5, 28)    <= sub_wire3(28);
	sub_wire1(5, 29)    <= sub_wire3(29);
	sub_wire1(5, 30)    <= sub_wire3(30);
	sub_wire1(5, 31)    <= sub_wire3(31);
	sub_wire1(4, 0)    <= sub_wire4(0);
	sub_wire1(4, 1)    <= sub_wire4(1);
	sub_wire1(4, 2)    <= sub_wire4(2);
	sub_wire1(4, 3)    <= sub_wire4(3);
	sub_wire1(4, 4)    <= sub_wire4(4);
	sub_wire1(4, 5)    <= sub_wire4(5);
	sub_wire1(4, 6)    <= sub_wire4(6);
	sub_wire1(4, 7)    <= sub_wire4(7);
	sub_wire1(4, 8)    <= sub_wire4(8);
	sub_wire1(4, 9)    <= sub_wire4(9);
	sub_wire1(4, 10)    <= sub_wire4(10);
	sub_wire1(4, 11)    <= sub_wire4(11);
	sub_wire1(4, 12)    <= sub_wire4(12);
	sub_wire1(4, 13)    <= sub_wire4(13);
	sub_wire1(4, 14)    <= sub_wire4(14);
	sub_wire1(4, 15)    <= sub_wire4(15);
	sub_wire1(4, 16)    <= sub_wire4(16);
	sub_wire1(4, 17)    <= sub_wire4(17);
	sub_wire1(4, 18)    <= sub_wire4(18);
	sub_wire1(4, 19)    <= sub_wire4(19);
	sub_wire1(4, 20)    <= sub_wire4(20);
	sub_wire1(4, 21)    <= sub_wire4(21);
	sub_wire1(4, 22)    <= sub_wire4(22);
	sub_wire1(4, 23)    <= sub_wire4(23);
	sub_wire1(4, 24)    <= sub_wire4(24);
	sub_wire1(4, 25)    <= sub_wire4(25);
	sub_wire1(4, 26)    <= sub_wire4(26);
	sub_wire1(4, 27)    <= sub_wire4(27);
	sub_wire1(4, 28)    <= sub_wire4(28);
	sub_wire1(4, 29)    <= sub_wire4(29);
	sub_wire1(4, 30)    <= sub_wire4(30);
	sub_wire1(4, 31)    <= sub_wire4(31);
	sub_wire1(3, 0)    <= sub_wire5(0);
	sub_wire1(3, 1)    <= sub_wire5(1);
	sub_wire1(3, 2)    <= sub_wire5(2);
	sub_wire1(3, 3)    <= sub_wire5(3);
	sub_wire1(3, 4)    <= sub_wire5(4);
	sub_wire1(3, 5)    <= sub_wire5(5);
	sub_wire1(3, 6)    <= sub_wire5(6);
	sub_wire1(3, 7)    <= sub_wire5(7);
	sub_wire1(3, 8)    <= sub_wire5(8);
	sub_wire1(3, 9)    <= sub_wire5(9);
	sub_wire1(3, 10)    <= sub_wire5(10);
	sub_wire1(3, 11)    <= sub_wire5(11);
	sub_wire1(3, 12)    <= sub_wire5(12);
	sub_wire1(3, 13)    <= sub_wire5(13);
	sub_wire1(3, 14)    <= sub_wire5(14);
	sub_wire1(3, 15)    <= sub_wire5(15);
	sub_wire1(3, 16)    <= sub_wire5(16);
	sub_wire1(3, 17)    <= sub_wire5(17);
	sub_wire1(3, 18)    <= sub_wire5(18);
	sub_wire1(3, 19)    <= sub_wire5(19);
	sub_wire1(3, 20)    <= sub_wire5(20);
	sub_wire1(3, 21)    <= sub_wire5(21);
	sub_wire1(3, 22)    <= sub_wire5(22);
	sub_wire1(3, 23)    <= sub_wire5(23);
	sub_wire1(3, 24)    <= sub_wire5(24);
	sub_wire1(3, 25)    <= sub_wire5(25);
	sub_wire1(3, 26)    <= sub_wire5(26);
	sub_wire1(3, 27)    <= sub_wire5(27);
	sub_wire1(3, 28)    <= sub_wire5(28);
	sub_wire1(3, 29)    <= sub_wire5(29);
	sub_wire1(3, 30)    <= sub_wire5(30);
	sub_wire1(3, 31)    <= sub_wire5(31);
	sub_wire1(2, 0)    <= sub_wire6(0);
	sub_wire1(2, 1)    <= sub_wire6(1);
	sub_wire1(2, 2)    <= sub_wire6(2);
	sub_wire1(2, 3)    <= sub_wire6(3);
	sub_wire1(2, 4)    <= sub_wire6(4);
	sub_wire1(2, 5)    <= sub_wire6(5);
	sub_wire1(2, 6)    <= sub_wire6(6);
	sub_wire1(2, 7)    <= sub_wire6(7);
	sub_wire1(2, 8)    <= sub_wire6(8);
	sub_wire1(2, 9)    <= sub_wire6(9);
	sub_wire1(2, 10)    <= sub_wire6(10);
	sub_wire1(2, 11)    <= sub_wire6(11);
	sub_wire1(2, 12)    <= sub_wire6(12);
	sub_wire1(2, 13)    <= sub_wire6(13);
	sub_wire1(2, 14)    <= sub_wire6(14);
	sub_wire1(2, 15)    <= sub_wire6(15);
	sub_wire1(2, 16)    <= sub_wire6(16);
	sub_wire1(2, 17)    <= sub_wire6(17);
	sub_wire1(2, 18)    <= sub_wire6(18);
	sub_wire1(2, 19)    <= sub_wire6(19);
	sub_wire1(2, 20)    <= sub_wire6(20);
	sub_wire1(2, 21)    <= sub_wire6(21);
	sub_wire1(2, 22)    <= sub_wire6(22);
	sub_wire1(2, 23)    <= sub_wire6(23);
	sub_wire1(2, 24)    <= sub_wire6(24);
	sub_wire1(2, 25)    <= sub_wire6(25);
	sub_wire1(2, 26)    <= sub_wire6(26);
	sub_wire1(2, 27)    <= sub_wire6(27);
	sub_wire1(2, 28)    <= sub_wire6(28);
	sub_wire1(2, 29)    <= sub_wire6(29);
	sub_wire1(2, 30)    <= sub_wire6(30);
	sub_wire1(2, 31)    <= sub_wire6(31);
	sub_wire1(1, 0)    <= sub_wire7(0);
	sub_wire1(1, 1)    <= sub_wire7(1);
	sub_wire1(1, 2)    <= sub_wire7(2);
	sub_wire1(1, 3)    <= sub_wire7(3);
	sub_wire1(1, 4)    <= sub_wire7(4);
	sub_wire1(1, 5)    <= sub_wire7(5);
	sub_wire1(1, 6)    <= sub_wire7(6);
	sub_wire1(1, 7)    <= sub_wire7(7);
	sub_wire1(1, 8)    <= sub_wire7(8);
	sub_wire1(1, 9)    <= sub_wire7(9);
	sub_wire1(1, 10)    <= sub_wire7(10);
	sub_wire1(1, 11)    <= sub_wire7(11);
	sub_wire1(1, 12)    <= sub_wire7(12);
	sub_wire1(1, 13)    <= sub_wire7(13);
	sub_wire1(1, 14)    <= sub_wire7(14);
	sub_wire1(1, 15)    <= sub_wire7(15);
	sub_wire1(1, 16)    <= sub_wire7(16);
	sub_wire1(1, 17)    <= sub_wire7(17);
	sub_wire1(1, 18)    <= sub_wire7(18);
	sub_wire1(1, 19)    <= sub_wire7(19);
	sub_wire1(1, 20)    <= sub_wire7(20);
	sub_wire1(1, 21)    <= sub_wire7(21);
	sub_wire1(1, 22)    <= sub_wire7(22);
	sub_wire1(1, 23)    <= sub_wire7(23);
	sub_wire1(1, 24)    <= sub_wire7(24);
	sub_wire1(1, 25)    <= sub_wire7(25);
	sub_wire1(1, 26)    <= sub_wire7(26);
	sub_wire1(1, 27)    <= sub_wire7(27);
	sub_wire1(1, 28)    <= sub_wire7(28);
	sub_wire1(1, 29)    <= sub_wire7(29);
	sub_wire1(1, 30)    <= sub_wire7(30);
	sub_wire1(1, 31)    <= sub_wire7(31);
	sub_wire1(0, 0)    <= sub_wire8(0);
	sub_wire1(0, 1)    <= sub_wire8(1);
	sub_wire1(0, 2)    <= sub_wire8(2);
	sub_wire1(0, 3)    <= sub_wire8(3);
	sub_wire1(0, 4)    <= sub_wire8(4);
	sub_wire1(0, 5)    <= sub_wire8(5);
	sub_wire1(0, 6)    <= sub_wire8(6);
	sub_wire1(0, 7)    <= sub_wire8(7);
	sub_wire1(0, 8)    <= sub_wire8(8);
	sub_wire1(0, 9)    <= sub_wire8(9);
	sub_wire1(0, 10)    <= sub_wire8(10);
	sub_wire1(0, 11)    <= sub_wire8(11);
	sub_wire1(0, 12)    <= sub_wire8(12);
	sub_wire1(0, 13)    <= sub_wire8(13);
	sub_wire1(0, 14)    <= sub_wire8(14);
	sub_wire1(0, 15)    <= sub_wire8(15);
	sub_wire1(0, 16)    <= sub_wire8(16);
	sub_wire1(0, 17)    <= sub_wire8(17);
	sub_wire1(0, 18)    <= sub_wire8(18);
	sub_wire1(0, 19)    <= sub_wire8(19);
	sub_wire1(0, 20)    <= sub_wire8(20);
	sub_wire1(0, 21)    <= sub_wire8(21);
	sub_wire1(0, 22)    <= sub_wire8(22);
	sub_wire1(0, 23)    <= sub_wire8(23);
	sub_wire1(0, 24)    <= sub_wire8(24);
	sub_wire1(0, 25)    <= sub_wire8(25);
	sub_wire1(0, 26)    <= sub_wire8(26);
	sub_wire1(0, 27)    <= sub_wire8(27);
	sub_wire1(0, 28)    <= sub_wire8(28);
	sub_wire1(0, 29)    <= sub_wire8(29);
	sub_wire1(0, 30)    <= sub_wire8(30);
	sub_wire1(0, 31)    <= sub_wire8(31);
	result    <= sub_wire9(31 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 8,
		lpm_type => "LPM_MUX",
		lpm_width => 32,
		lpm_widths => 3
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire9
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
-- Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
-- Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
-- Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
-- Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
-- Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
-- Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL "sel[2..0]"
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 2 32 0 data2x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 3 32 0 data3x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 4 32 0 data4x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 5 32 0 data5x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 6 32 0 data6x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 7 32 0 data7x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux3to8_32bit.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux3to8_32bit.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux3to8_32bit.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux3to8_32bit.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux3to8_32bit_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
