MUX1TO2_29BIT_inst : MUX1TO2_29BIT PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
