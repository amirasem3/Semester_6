LAND_inst : LAND PORT MAP (
		result	 => result_sig
	);
