ISUB_inst : ISUB PORT MAP (
		result	 => result_sig
	);
