lADD_inst : lADD PORT MAP (
		result	 => result_sig
	);
