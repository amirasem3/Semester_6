retn_inst : retn PORT MAP (
		result	 => result_sig
	);
