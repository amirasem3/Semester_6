AORB_inst : AORB PORT MAP (
		result	 => result_sig
	);
