module rom(address,data);
input [6:0] address; //needs to be changed
output [22:0] data;	//needs to be changed
reg [22:0] array[126:0];	//needs to be changed
always @*
begin
array[0] = 23'b00010001000000001011011;              //fetch
array[1] = 23'b00000000000000000000000;              //nop
array[2] = 23'b01000010000100000000011;              //BIPUSH
array[3] = 23'b00000001001000000000000;              //
array[4] = 23'b00000000001100000000000;              //GOTO
array[5] = 23'b00100011000000000000110;              //IADD
array[6] = 23'b00000000000000000000111;              //
array[7] = 23'b00000000010100000001000;              //
array[8] = 23'b00000100000000000000000;              //
array[9] = 23'b00100011000000000001010;              //IFEQ
array[10] = 23'b00000000000011000001100;              //
array[11] = 23'b00000000001100000001100;              //
array[12] = 23'b00000001000000000001101;              //
array[13] = 23'b00000001000000000000000;              //
array[14] = 23'b00100011000000000001111;              //IFLT
array[15] = 23'b00000000000001000010010;              //
array[16] = 23'b00000001000000000010001;              //
array[17] = 23'b00000001000000000000000;              //
array[18] = 23'b00000000001100000000000;              //
array[19] = 23'b00100011000000000010100;              //If_icmpeq
array[20] = 23'b00110011000000000010101;              //
array[21] = 23'b00000000010000000010110;              //
array[22] = 23'b00000000100000000010111;              //
array[23] = 23'b00000000000010000011001;              //
array[24] = 23'b00000000001100000000000;              //
array[25] = 23'b00000001000000000011010;              //
array[26] = 23'b00000001000000000000000;              //
array[27] = 23'b01000000000100000011100;              //Iinc
array[28] = 23'b01010001000000000011101;              //
array[29] = 23'b10010000000000000011110;              //
array[30] = 23'b01000001000100000011111;              //
array[31] = 23'b00000000100100000100000;              //
array[32] = 23'b00000000010100000100001;              //
array[33] = 23'b00000101000000000000000;              //
array[34] = 23'b01000000000100000100011;              //ILOAD
array[35] = 23'b01010001000000000100100;              //
array[36] = 23'b10010010000000000100101;              //
array[37] = 23'b00000000011100000000000;              //
array[38] = 23'b00100011000000000100111;              //IStore
array[39] = 23'b01000000000000000101000;              //
array[40] = 23'b00000000000100000101001;              //
array[41] = 23'b01010001000000000101010;              //
array[42] = 23'b00001000000000000000000;              //
array[43] = 23'b00100011000000000101100;              //ISUB
array[44] = 23'b00110000000000000101101;              //
array[45] = 23'b00000000010000000101110;              //
array[46] = 23'b00000100000000000000000;              //
array[47] = 23'b00100010000000000110000;              //DUP
array[48] = 23'b00000000011100000000000;              //
array[49] = 23'b00100011000000000110010;              //LAND
array[50] = 23'b00110000000000000110011;              //
array[51] = 23'b01110000000000000110100;              //
array[52] = 23'b00000100000000000000000;              //
array[53] = 23'b00100011000000000110110;              //swap
array[54] = 23'b00110000000000000110111;              //
array[55] = 23'b00000010011100000111000;              //
array[56] = 23'b00000111000000000111001;              //
array[57] = 23'b00000100000000000000000;              //
array[58] = 23'b10110000000000000000000;              //wide
array[59] = 23'b00100011000000000111100;              //IOR
array[60] = 23'b00110000000000000111101;              //
array[61] = 23'b10000000000000000111110;              //
array[62] = 23'b00000100000000000000000;              //
array[63] = 23'b00000000101100001000000;              //LDC_W
array[64] = 23'b00000010101000001000001;              //
array[65] = 23'b00000000011100000000000;              //
array[66] = 23'b00000011000000000000000;              //POP
array[67] = 23'b10100001000000001000100;              //LDASP
array[68] = 23'b00000001000000001000101;              //
array[69] = 23'b00000001000000001000110;              //
array[70] = 23'b00000001000000000000000;              //
array[71] = 23'b01101010000000001001000;              //ENVOKE
array[72] = 23'b00001001000000001001001;              //
array[73] = 23'b11010001110000001001010;              //
array[74] = 23'b00000000100100001001011;              //
array[75] = 23'b00001011110100001001100;              //
array[76] = 23'b00001110000000001001101;              //
array[77] = 23'b00000000010000001001110;              //
array[78] = 23'b00000001111000001001111;              //
array[79] = 23'b00000000110000001010000;              //
array[80] = 23'b00000001100100001010001;              //
array[81] = 23'b00001011110100001010010;              //
array[82] = 23'b00001110000000001010011;              //
array[83] = 23'b00000001010100001010100;              //
array[84] = 23'b00001100000000001010101;              //
array[85] = 23'b00000010111100001010110;              //
array[86] = 23'b00001101000000000000000;              //
array[87] = 23'b00001010000000001011000;              //RETURN

array[88] = 23'b11110011000000001011001;              //
array[89] = 23'b00000000011000001011010;              //



array[90] = 23'b00001111000000000000000;              //
array[91] = 23'b00000000000000110000000;              
end
assign data=array[address];
endmodule