ISTORE_inst : ISTORE PORT MAP (
		result	 => result_sig
	);
