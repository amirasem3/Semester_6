BMA_inst : BMA PORT MAP (
		result	 => result_sig
	);
