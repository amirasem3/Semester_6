FETCH_inst : FETCH PORT MAP (
		result	 => result_sig
	);
