TESTCONSTANT_inst : TESTCONSTANT PORT MAP (
		result	 => result_sig
	);
