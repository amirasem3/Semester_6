ILOAD_inst : ILOAD PORT MAP (
		result	 => result_sig
	);
