AN_inst : AN PORT MAP (
		result	 => result_sig
	);
