LDASP_inst : LDASP PORT MAP (
		result	 => result_sig
	);
