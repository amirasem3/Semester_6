SHIF4L_inst : SHIF4L PORT MAP (
		result	 => result_sig
	);
