AANDB_inst : AANDB PORT MAP (
		result	 => result_sig
	);
