SWAP_inst : SWAP PORT MAP (
		result	 => result_sig
	);
