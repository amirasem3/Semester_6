BPA_inst : BPA PORT MAP (
		result	 => result_sig
	);
