IINC_inst : IINC PORT MAP (
		result	 => result_sig
	);
