A_inst : A PORT MAP (
		result	 => result_sig
	);
