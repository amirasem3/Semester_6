ENVOKE_inst : ENVOKE PORT MAP (
		result	 => result_sig
	);
