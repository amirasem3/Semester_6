IFLT_inst : IFLT PORT MAP (
		result	 => result_sig
	);
