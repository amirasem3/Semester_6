ZERO_inst : ZERO PORT MAP (
		result	 => result_sig
	);
