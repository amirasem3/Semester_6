POP_inst : POP PORT MAP (
		result	 => result_sig
	);
