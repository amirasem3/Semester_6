IFEQ_inst : IFEQ PORT MAP (
		result	 => result_sig
	);
